----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:46:09 10/05/2022 
-- Design Name: 
-- Module Name:    DBUF_reg8_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DBUF_reg8_1 is
    Port ( I_clk : in  STD_LOGIC;
           I_en : in  STD_LOGIC;
			  I_dir : in STD_LOGIC;
           I_data_buff : in  STD_LOGIC_VECTOR (7 downto 0);
           I_data_uct : in  STD_LOGIC_VECTOR (7 downto 0);
			  O_data_buff : out  STD_LOGIC_VECTOR (7 downto 0);
           O_data_uct : out  STD_LOGIC_VECTOR (7 downto 0));
end DBUF_reg8_1;

architecture Behavioral of DBUF_reg8_1 is

begin
	process(I_clk, I_en)
	begin
		if rising_edge(I_clk) and I_en='1' then
			if I_dir = '1' then
				O_data_uct <= I_data_buff;
			else
				O_data_buff <= I_data_uct;
			end if;
		end if;
	end process;

end Behavioral;

